module design1(iCLOCK, inRESET, iRESET_SYNC, iCTRL_HOLD, iPFLAGR_VALID, iPFLAGR, iPREV_INST_VALID, iPREV_BUSY, iPREV_FLAG_WRITE, iSHIFT_VALID, iSHIFT_FLAG, iADDER_VALID, iADDER_FLAG, iMUL_VALID, iMUL_FLAG, iLOGIC_VALID, iLOGIC_FLAG, oFLAG);
  wire [4:0] _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire [4:0] _04_;
  wire [4:0] _05_;
  wire [4:0] _06_;
  wire [4:0] _07_;
  wire [4:0] _08_;
  wire [4:0] _09_;
  wire [4:0] _10_;
  wire [4:0] _11_;
  wire [4:0] _12_;
  reg [4:0] b_sysreg_flags = 5'd0;
  input [4:0] iADDER_FLAG;
  input iADDER_VALID;
  input iCLOCK;
  input iCTRL_HOLD;
  input [4:0] iLOGIC_FLAG;
  input iLOGIC_VALID;
  input [4:0] iMUL_FLAG;
  input iMUL_VALID;
  input [4:0] iPFLAGR;
  input iPFLAGR_VALID;
  input iPREV_BUSY;
  input iPREV_FLAG_WRITE;
  input iPREV_INST_VALID;
  input iRESET_SYNC;
  input [4:0] iSHIFT_FLAG;
  input iSHIFT_VALID;
  input inRESET;
  output [4:0] oFLAG;
  assign _01_ = _02_ &&  iPREV_INST_VALID;
  assign _02_ = !  iPREV_BUSY;
  assign _03_ = !  inRESET;
  always @(posedge iCLOCK)
      b_sysreg_flags <= _00_;
  assign _04_ = iADDER_VALID ?  iADDER_FLAG : _12_;
  assign _05_ = iSHIFT_VALID ?  iSHIFT_FLAG : _04_;
  assign _06_ = iPREV_FLAG_WRITE ?  _05_ : b_sysreg_flags;
  assign _07_ = _01_ ?  _06_ : b_sysreg_flags;
  assign _08_ = iCTRL_HOLD ?  b_sysreg_flags : _07_;
  assign _09_ = iPFLAGR_VALID ?  iPFLAGR : _08_;
  assign _10_ = iRESET_SYNC ?  5'h00 : _09_;
  assign _00_ = _03_ ?  5'h00 : _10_;
  assign _11_ = iLOGIC_VALID ?  iLOGIC_FLAG : b_sysreg_flags;
  assign _12_ = iMUL_VALID ?  iMUL_FLAG : _11_;
  assign oFLAG = b_sysreg_flags;
endmodule

module design2(iLOGIC_VALID, iPFLAGR, iSHIFT_FLAG, iMUL_FLAG, iSHIFT_VALID, iADDER_FLAG, inRESET, iLOGIC_FLAG, iADDER_VALID, iPFLAGR_VALID, iPREV_FLAG_WRITE, iPREV_INST_VALID, iMUL_VALID, iCTRL_HOLD, iRESET_SYNC, iPREV_BUSY, iCLOCK, oFLAG);
input  iLOGIC_VALID;
input [4:0] iPFLAGR;
input [4:0] iSHIFT_FLAG;
input [4:0] iMUL_FLAG;
input  iSHIFT_VALID;
input [4:0] iADDER_FLAG;
input  inRESET;
input [4:0] iLOGIC_FLAG;
input  iADDER_VALID;
input  iPFLAGR_VALID;
input  iPREV_FLAG_WRITE;
input  iPREV_INST_VALID;
input  iMUL_VALID;
input  iCTRL_HOLD;
input  iRESET_SYNC;
input  iPREV_BUSY;
input  iCLOCK;
output [4:0] oFLAG;
reg [4:0] b_sysreg_flags = 5'd0;
wire  _01_;
wire [4:0] _11_;
wire [4:0] _05_;
wire [4:0] _04_;
wire  _02_;
wire [4:0] _09_;
wire [4:0] _10_;
wire [4:0] _06_;
wire [4:0] _08_;
wire [4:0] _00_;
wire  _03_;
wire [4:0] _12_;
wire [4:0] _07_;
always @(posedge iCLOCK)
    b_sysreg_flags <= _00_;
assign _01_ = (_02_) && (iPREV_INST_VALID);
assign _11_ = (iLOGIC_VALID) ? (iLOGIC_FLAG) : (b_sysreg_flags);
assign _05_ = (iSHIFT_VALID) ? (iSHIFT_FLAG) : (_04_);
assign _04_ = (iADDER_VALID) ? (iADDER_FLAG) : (_12_);
assign _02_ = !(iPREV_BUSY);
assign _09_ = (iPFLAGR_VALID) ? (iPFLAGR) : (_08_);
assign _10_ = (iRESET_SYNC) ? (5'h0) : (_09_);
assign _06_ = (iPREV_FLAG_WRITE) ? (_05_) : (b_sysreg_flags);
assign _08_ = (iCTRL_HOLD) ? (b_sysreg_flags) : (_07_);
assign _00_ = (_03_) ? (5'h0) : (_10_);
assign _03_ = !(inRESET);
assign _12_ = (iMUL_VALID) ? (iMUL_FLAG) : (_11_);
assign _07_ = (_01_) ? (_06_) : (b_sysreg_flags);
assign oFLAG = b_sysreg_flags;
endmodule

module miter();
wire [4:0] oFLAG1, oFLAG2;
design1 inst1 (.iCLOCK(iCLOCK),.inRESET(inRESET),.iRESET_SYNC(iRESET_SYNC),.iCTRL_HOLD(iCTRL_HOLD),.iPFLAGR_VALID(iPFLAGR_VALID),.iPFLAGR(iPFLAGR),.iPREV_INST_VALID(iPREV_INST_VALID),.iPREV_BUSY(iPREV_BUSY),.iPREV_FLAG_WRITE(iPREV_FLAG_WRITE),.iSHIFT_VALID(iSHIFT_VALID),.iSHIFT_FLAG(iSHIFT_FLAG),.iADDER_VALID(iADDER_VALID),.iADDER_FLAG(iADDER_FLAG),.iMUL_VALID(iMUL_VALID),.iMUL_FLAG(iMUL_FLAG),.iLOGIC_VALID(iLOGIC_VALID),.iLOGIC_FLAG(iLOGIC_FLAG),.oFLAG(oFLAG1));
design2 inst2 (.iCLOCK(iCLOCK),.inRESET(inRESET),.iRESET_SYNC(iRESET_SYNC),.iCTRL_HOLD(iCTRL_HOLD),.iPFLAGR_VALID(iPFLAGR_VALID),.iPFLAGR(iPFLAGR),.iPREV_INST_VALID(iPREV_INST_VALID),.iPREV_BUSY(iPREV_BUSY),.iPREV_FLAG_WRITE(iPREV_FLAG_WRITE),.iSHIFT_VALID(iSHIFT_VALID),.iSHIFT_FLAG(iSHIFT_FLAG),.iADDER_VALID(iADDER_VALID),.iADDER_FLAG(iADDER_FLAG),.iMUL_VALID(iMUL_VALID),.iMUL_FLAG(iMUL_FLAG),.iLOGIC_VALID(iLOGIC_VALID),.iLOGIC_FLAG(iLOGIC_FLAG),.oFLAG(oFLAG2));
always @(posedge clk) begin
assert(oFLAG1 == oFLAG2);
end
endmodule