module module_6(rc_reqn, rstn, rc_is_idle, clk, rc_ackn);
input  rc_reqn;
input  rstn;
input  rc_is_idle;
input  clk;
output  rc_ackn;
reg [1:0] state_c;
wire  _11_;
wire  _10_;
wire  _01_;
wire [1:0] _00_;
wire  _04_;
wire [1:0] state_n;
wire  _07_;
wire  _05_;
wire [1:0] _06_;
wire  _09_;
wire  _08_;
wire  _03_;
wire [1:0] _12_;
wire [1:0] _02_;
always @(posedge clk)
    state_c <= _00_;
assign _11_ = (rc_is_idle) ? (1'h0) : (1'h1);
assign _10_ = (state_c) == (2'h1);
assign _01_ = (_05_) ? (_11_) : (1'hx);
assign _00_ = (_04_) ? (2'h0) : (state_n);
assign _04_ = !(rstn);
assign state_n = (_09_ ? _12_ : (_08_ ? _02_ : 2'h0));
assign _07_ = (state_c) == (2'h1);
assign _05_ = (state_c) == (2'h1);
assign _06_ = (rc_is_idle) ? (2'h0) : (2'h1);
assign _09_ = (state_c) == (2'h0);
assign _08_ = (state_c) == (2'h1);
assign _03_ = !(rc_reqn);
assign _12_ = (_03_) ? (2'h1) : (2'h0);
assign _02_ = (_07_) ? (_06_) : (2'hx);
assign rc_ackn = (_10_) ? (_01_) : (1'h1);
endmodule