module vga_text(clk25mhz, hindex, vindex, standard, emphasized, background, char_data, font_data, char_address, font_address, color);
  wire [2:0] _00_;
  wire [11:0] _01_;
  wire [2:0] _02_;
  wire [3:0] _03_;
  wire [2:0] _04_;
  wire [3:0] _05_;
  wire [31:0] _06_;
  wire [31:0] _07_;
  wire [31:0] _08_;
  wire _09_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire _15_;
  wire _16_;
  wire _17_;
  wire _18_;
  wire _19_;
  wire _20_;
  wire _21_;
  wire _22_;
  wire _23_;
  wire _24_;
  wire _25_;
  wire [2:0] _26_;
  wire [2:0] _27_;
  wire [3:0] _28_;
  wire [3:0] _29_;
  wire [3:0] _30_;
  wire [2:0] _31_;
  wire [2:0] _32_;
  wire [11:0] _33_;
  wire [11:0] _34_;
  wire [11:0] _35_;
  wire [11:0] _36_;
  wire [11:0] _37_;
  wire _38_;
  wire [31:0] _39_;
  input [3:0] background;
  reg [2:0] bright = 3'h0;
  output [11:0] char_address;
  reg [11:0] char_address = 12'h000;
  reg [2:0] char_col = 3'h0;
  input [7:0] char_data;
  reg [3:0] char_row = 4'h0;
  input clk25mhz;
  output [7:0] color;
  reg [2:0] dark = 3'h0;
  input [3:0] emphasized;
  output [9:0] font_address;
  reg [9:0] font_address;
  input [13:0] font_data;
  reg [3:0] foreground;
  input [9:0] hindex;
  wire [3:0] pixel_color;
  input [3:0] standard;
  input [9:0] vindex;
  assign _06_ = char_address +  32'd1;
  assign _07_ = char_col +  32'd1;
  assign _08_ = char_row +  32'd1;
  assign _09_ = _38_ ==  32'd1;
  assign _10_ = char_col ==  32'd7;
  assign _11_ = hindex ==  32'd640;
  assign _12_ = char_row ==  32'd13;
  assign _13_ = char_address ==  32'd2720;
  assign _14_ = char_data[7] ==  32'd1;
  assign _15_ = pixel_color[3] ==  32'd1;
  assign _16_ = pixel_color[2:0] ==  32'd0;
  assign _17_ = vindex >=  32'd2;
  assign _18_ = hindex >  32'd0;
  assign _19_ = _17_ &&  _22_;
  assign _20_ = _18_ &&  _24_;
  assign _21_ = _20_ &&  _25_;
  assign _22_ = vindex <  32'd478;
  assign _23_ = hindex <  32'd640;
  assign _24_ = hindex <  32'd641;
  assign _25_ = vindex <  32'd480;
  always @(posedge clk25mhz)
      dark <= _04_;
  always @(posedge clk25mhz)
      bright <= _00_;
  always @(posedge clk25mhz)
      font_address <= { char_data[6:0], char_col };
  always @(posedge clk25mhz)
      foreground <= _05_;
  always @(posedge clk25mhz)
      char_address <= _01_;
  always @(posedge clk25mhz)
      char_col <= _02_;
  always @(posedge clk25mhz)
      char_row <= _03_;
  assign _26_ = _16_ ?  3'h7 : pixel_color[2:0];
  assign _27_ = _15_ ?  _26_ : 3'h0;
  assign _00_ = _21_ ?  _27_ : 3'h0;
  assign _04_ = _21_ ?  pixel_color[2:0] : 3'h0;
  assign _28_ = _12_ ?  4'h0 : _08_[3:0];
  assign _29_ = _11_ ?  _28_ : char_row;
  assign _30_ = _23_ ?  char_row : _29_;
  assign _03_ = _19_ ?  _30_ : char_row;
  assign _31_ = _10_ ?  3'h0 : _07_[2:0];
  assign _32_ = _23_ ?  _31_ : char_col;
  assign _02_ = _19_ ?  _32_ : char_col;
  assign _33_ = _13_ ?  12'h000 : char_address;
  assign _34_ = _12_ ?  _33_ : _39_[11:0];
  assign _35_ = _11_ ?  _34_ : char_address;
  assign _36_ = _10_ ?  _06_[11:0] : char_address;
  assign _37_ = _23_ ?  _36_ : _35_;
  assign _01_ = _19_ ?  _37_ : char_address;
  wire [13:0] _88_ = font_data;
  assign _38_ = _88_[char_row +: 1];
  assign _39_ = char_address -  32'd80;
  assign pixel_color = _09_ ?  foreground : background;
  assign _05_ = _14_ ?  emphasized : standard;
  assign color = { dark[2], bright[2], 1'h0, dark[1], bright[1], 1'h0, dark[0], bright[0] };
endmodule