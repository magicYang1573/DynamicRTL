module module_8(we, reset_in, addr, mclk28, bank1, card_ram_we, card_ram_rd, ram_addr);
input  we;
input  reset_in;
input [15:0] addr;
input  mclk28;
output  bank1;
output  card_ram_we;
output  card_ram_rd;
output [17:0] ram_addr;
reg  bank1;
reg  pre_wr_en;
reg  bankB;
reg  sat_write_en;
reg  write_en;
reg  sat_pre_wr_en;
reg [2:0] bank16k;
reg  read_en;
reg  sat_read_en;
reg [15:0] addr2;
wire  _001_;
wire  _047_;
wire  _012_;
wire  _027_;
wire  _029_;
wire  _013_;
wire  _003_;
wire  _021_;
wire  _033_;
wire [2:0] _000_;
wire  _016_;
wire  _022_;
wire  _045_;
wire  Dxxx;
wire  _028_;
wire  _004_;
wire  _018_;
wire  _048_;
wire  _019_;
wire  _043_;
wire  _002_;
wire  _039_;
wire  _017_;
wire  _031_;
wire  _014_;
wire  _038_;
wire  _023_;
wire  _007_;
wire  _025_;
wire  _037_;
wire  _009_;
wire  _040_;
wire  _011_;
wire  _036_;
wire  _049_;
wire  _010_;
wire [2:0] _034_;
wire  _042_;
wire  _020_;
wire  _030_;
wire  _041_;
wire  _024_;
wire  _032_;
wire  _006_;
wire  _005_;
wire  _046_;
wire  _015_;
wire [2:0] _035_;
wire  DEF;
wire  _026_;
wire  _008_;
wire  _044_;
always @(posedge mclk28)
    bank1 <= _001_;
always @(posedge mclk28)
    pre_wr_en <= _003_;
always @(posedge mclk28)
    bankB <= _002_;
always @(posedge mclk28)
    sat_write_en <= _007_;
always @(posedge mclk28)
    write_en <= _008_;
always @(posedge mclk28)
    sat_pre_wr_en <= _005_;
always @(posedge mclk28)
    bank16k <= _000_;
always @(posedge mclk28)
    read_en <= _004_;
always @(posedge mclk28)
    sat_read_en <= _006_;
always @(posedge mclk28)
    addr2 <= addr;
assign _001_ = (reset_in) ? (1'h0) : (_047_);
assign _047_ = (_009_) ? (addr[3:3]) : (bank1);
assign _012_ = (_011_) & (_029_);
assign _027_ = (addr[13:12]) != (2'h0);
assign _029_ = !(we);
assign _013_ = (_020_) & (_026_);
assign _003_ = (reset_in) ? (1'h0) : (_044_);
assign _021_ = (addr[2:2]) == (32'd0);
assign _033_ = !(_017_);
assign _000_ = (reset_in) ? (bank16k) : (_035_);
assign _016_ = (addr[12:12]) & (_032_);
assign _022_ = (addr[15:14]) == (2'h3);
assign _045_ = (_009_) ? (_012_) : (write_en);
assign Dxxx = (addr[15:12]) == (4'hd);
assign _028_ = !(we);
assign _004_ = (reset_in) ? (1'h0) : (_046_);
assign _018_ = (addr[12:12]) & (_033_);
assign _048_ = (addr[0:0]) ^ (addr[1:1]);
assign _019_ = (addr[15:4]) == (32'd3080);
assign _043_ = (_013_) ? (_042_) : (bankB);
assign _002_ = (reset_in) ? (1'h0) : (_043_);
assign _039_ = (_013_) ? (_038_) : (sat_write_en);
assign _017_ = (bank1) & (Dxxx);
assign _031_ = !(_049_);
assign _014_ = (addr[0:0]) & (sat_pre_wr_en);
assign _038_ = (_021_) ? (_014_) : (sat_write_en);
assign _023_ = (_024_) && (DEF);
assign _007_ = (reset_in) ? (1'h0) : (_039_);
assign _025_ = (addr2) != (addr);
assign _037_ = (_013_) ? (_036_) : (sat_pre_wr_en);
assign _009_ = (_019_) & (_025_);
assign _040_ = (_021_) ? (_031_) : (sat_read_en);
assign _011_ = (addr[0:0]) & (pre_wr_en);
assign _036_ = (_021_) ? (addr[0:0]) : (sat_pre_wr_en);
assign _049_ = (addr[0:0]) ^ (addr[1:1]);
assign _010_ = (addr[0:0]) & (_028_);
assign _034_ = (_021_) ? (bank16k) : ({addr[3:3], addr[1:0]});
assign _042_ = (_021_) ? (addr[3:3]) : (bankB);
assign _020_ = (addr[15:4]) == (32'd3085);
assign _030_ = !(_048_);
assign _041_ = (_013_) ? (_040_) : (sat_read_en);
assign _024_ = (sat_write_en) || (sat_read_en);
assign _032_ = !(_015_);
assign _006_ = (reset_in) ? (1'h0) : (_041_);
assign _005_ = (reset_in) ? (1'h0) : (_037_);
assign _046_ = (_009_) ? (_030_) : (read_en);
assign _015_ = (bankB) & (Dxxx);
assign _035_ = (_013_) ? (_034_) : (bank16k);
assign DEF = (_022_) & (_027_);
assign _026_ = (addr2) != (addr);
assign _008_ = (reset_in) ? (1'h1) : (_045_);
assign _044_ = (_009_) ? (_010_) : (pre_wr_en);
assign card_ram_we = (write_en) | (sat_write_en);
assign card_ram_rd = (read_en) | (sat_read_en);
assign ram_addr = (_023_) ? ({1'h1, bank16k, addr[13:13], _016_, addr[11:0]}) : ({2'h0, addr[15:13], _018_, addr[11:0]});
endmodule